
import ClientServer ::*;
import Complex      ::*;
import FIFO         ::*;
import Reg6375      ::*;
import GetPut       ::*;
import Real         ::*;
import Vector       ::*;
import BRAMFIFO     ::*;

import AudioProcessorTypes::*;

typedef Server#(
    Vector#(FFT_POINTS, ComplexSample),
    Vector#(FFT_POINTS, ComplexSample)
) FFT;

// Get the appropriate twiddle factor for the given stage and index.
// This computes the twiddle factor statically.
function ComplexSample getTwiddle(Integer stage, Integer index, Integer points);
    Integer i = ((2*index)/(2 ** (log2(points)-stage))) * (2 ** (log2(points)-stage));
    return cmplx(fromReal(cos(fromInteger(i)*pi/fromInteger(points))),
                 fromReal(-1*sin(fromInteger(i)*pi/fromInteger(points))));
endfunction

// Generate a table of all the needed twiddle factors.
// The table can be used for looking up a twiddle factor dynamically.
typedef Vector#(FFT_LOG_POINTS, Vector#(TDiv#(FFT_POINTS, 2), ComplexSample)) TwiddleTable;
function TwiddleTable genTwiddles();
    TwiddleTable twids = newVector;
    for (Integer s = 0; s < valueof(FFT_LOG_POINTS); s = s+1) begin
        for (Integer i = 0; i < valueof(TDiv#(FFT_POINTS, 2)); i = i+1) begin
            twids[s][i] = getTwiddle(s, i, valueof(FFT_POINTS));
        end
    end
    return twids;
endfunction

// Given the destination location and the number of points in the fft, return
// the source index for the permutation.
function Integer permute(Integer dst, Integer points);
    Integer src = ?;
    if (dst < points/2) begin
        src = dst*2;
    end else begin
        src = (dst - points/2)*2 + 1;
    end
    return src;
endfunction

// Reorder the given vector by swapping words at positions
// corresponding to the bit-reversal of their indices.
// The reordering can be done either as as the
// first or last phase of the FFT transformation.
function Vector#(FFT_POINTS, ComplexSample) bitReverse(Vector#(FFT_POINTS,ComplexSample) inVector);
    Vector#(FFT_POINTS, ComplexSample) outVector = newVector();
    for(Integer i = 0; i < valueof(FFT_POINTS); i = i+1) begin
        Bit#(FFT_LOG_POINTS) reversal = reverseBits(fromInteger(i));
        outVector[reversal] = inVector[i];
    end
    return outVector;
endfunction

function Vector#(FFT_POINTS, ComplexSample) aebitReverse(Vector#(FFT_POINTS,ComplexSample) inVector);
  Vector#(FFT_POINTS, ComplexSample) outVector = newVector();
  // hardcoded for 8-pt fft.
  // for(Integer i = 0; i < valueof(FFT_POINTS); i = i+1) begin
  //     Bit#(FFT_LOG_POINTS) reversal = reverseBits(fromInteger(i));
  //     outVector[reversal] = inVector[i];
  // end
  outVector[0] = inVector[0];
  outVector[4] = inVector[1];
  outVector[2] = inVector[2];
  outVector[6] = inVector[3];
  outVector[1] = inVector[4];
  outVector[5] = inVector[5];
  outVector[3] = inVector[6];
  outVector[7] = inVector[7];
  return outVector;
endfunction

// 2-way Butterfly
function Vector#(2, ComplexSample) bfly2(Vector#(2, ComplexSample) t, ComplexSample k);
    ComplexSample m = t[1] * k;

    Vector#(2, ComplexSample) z = newVector();
    z[0] = t[0] + m;
    z[1] = t[0] - m;

    return z;
endfunction

// Perform a single stage of the FFT, consisting of butterflys and a single
// permutation.
// We pass the table of twiddles as an argument so we can look those up
// dynamically if need be.
function Vector#(FFT_POINTS, ComplexSample) stage_ft(TwiddleTable twiddles, Bit#(TLog#(FFT_LOG_POINTS)) stage, Vector#(FFT_POINTS, ComplexSample) stage_in);
    Vector#(FFT_POINTS, ComplexSample) stage_temp = newVector();
    for(Integer i = 0; i < (valueof(FFT_POINTS)/2); i = i+1) begin
        Integer idx = i * 2;
        let twid = twiddles[stage][i];
        let y = bfly2(takeAt(idx, stage_in), twid);

        stage_temp[idx]   = y[0];
        stage_temp[idx+1] = y[1];
    end

    Vector#(FFT_POINTS, ComplexSample) stage_out = newVector();
    for (Integer i = 0; i < valueof(FFT_POINTS); i = i+1) begin
        stage_out[i] = stage_temp[permute(i, valueof(FFT_POINTS))];
    end
    return stage_out;
endfunction

function Vector#(FFT_POINTS, ComplexSample) ae_stage_ft(TwiddleTable twiddles, Bit#(TLog#(FFT_LOG_POINTS)) stage, Vector#(FFT_POINTS, ComplexSample) stage_in);
  Vector#(FFT_POINTS, ComplexSample) stage_temp = newVector();
  // hard coded for 8-pt fft.
  // for(Integer i = 0; i < (valueof(FFT_POINTS)/2); i = i+1) begin
  //     Integer idx = i * 2;
  //     let twid = twiddles[stage][i];
  //     let y = bfly2(takeAt(idx, stage_in), twid);

  //     stage_temp[idx]   = y[0];
  //     stage_temp[idx+1] = y[1];
  // end
  let y0 = bfly2(takeAt(0, stage_in), twiddles[stage][0]);
  stage_temp[0] = y0[0];
  stage_temp[1] = y0[1];
  let y1 = bfly2(takeAt(2, stage_in), twiddles[stage][2]);
  stage_temp[2] = y1[0];
  stage_temp[3] = y1[1];
  let y2 = bfly2(takeAt(4, stage_in), twiddles[stage][4]);
  stage_temp[4] = y2[0];
  stage_temp[5] = y2[1];
  let y3 = bfly2(takeAt(6, stage_in), twiddles[stage][6]);
  stage_temp[6] = y3[0];
  stage_temp[7] = y3[1];

  Vector#(FFT_POINTS, ComplexSample) stage_out = newVector();
  // hardcoded for 8-pt fft.
  // for (Integer i = 0; i < valueof(FFT_POINTS); i = i+1) begin
  //     stage_out[i] = stage_temp[permute(i, valueof(FFT_POINTS))];
  // end
  stage_out[0] = stage_temp[0];
  stage_out[1] = stage_temp[4];
  stage_out[2] = stage_temp[1];
  stage_out[3] = stage_temp[5];
  stage_out[4] = stage_temp[2];
  stage_out[5] = stage_temp[6];
  stage_out[6] = stage_temp[3];
  stage_out[7] = stage_temp[7];
  return stage_out;
endfunction

module mkCombinationalFFT (FFT);

  // Statically generate the twiddle factors table.
  TwiddleTable twiddles = genTwiddles();

  // Define the stage_f function which uses the generated twiddles.
  function Vector#(FFT_POINTS, ComplexSample) stage_f(Bit#(TLog#(FFT_LOG_POINTS)) stage, Vector#(FFT_POINTS, ComplexSample) stage_in);
      return stage_ft(twiddles, stage, stage_in);
  endfunction

  FIFO#(Vector#(FFT_POINTS, ComplexSample)) inputFIFO  <- mkSizedBRAMFIFO(1);
  FIFO#(Vector#(FFT_POINTS, ComplexSample)) outputFIFO <- mkSizedBRAMFIFO(1);

  // This rule performs fft using a big mass of combinational logic.
  rule comb_fft;

    Vector#(TAdd#(1, FFT_LOG_POINTS), Vector#(FFT_POINTS, ComplexSample)) stage_data = newVector();
    stage_data[0] = inputFIFO.first();
    inputFIFO.deq();

    for(Integer stage = 0; stage < valueof(FFT_LOG_POINTS); stage=stage+1) begin
        stage_data[stage+1] = stage_f(fromInteger(stage), stage_data[stage]);
    end

    outputFIFO.enq(stage_data[valueof(FFT_LOG_POINTS)]);
  endrule

  interface Put request;
    method Action put(Vector#(FFT_POINTS, ComplexSample) x);
        inputFIFO.enq(bitReverse(x));
    endmethod
  endinterface

  interface Get response = toGet(outputFIFO);

endmodule

module mkPipelinedFFT (FFT);

  // Statically generate the twiddle factors table.
  TwiddleTable twiddles = genTwiddles();

  // Define the stage_f function which uses the generated twiddles.
  function Vector#(FFT_POINTS, ComplexSample) stage_f(Bit#(TLog#(FFT_LOG_POINTS)) stage, Vector#(FFT_POINTS, ComplexSample) stage_in);
      return stage_ft(twiddles, stage, stage_in);
  endfunction

  FIFO#(Vector#(FFT_POINTS, ComplexSample)) inputFIFO  <- mkSizedBRAMFIFO(1);
  FIFO#(Vector#(FFT_POINTS, ComplexSample)) isb1  <- mkSizedBRAMFIFO(1);
  FIFO#(Vector#(FFT_POINTS, ComplexSample)) isb2  <- mkSizedBRAMFIFO(1);
  FIFO#(Vector#(FFT_POINTS, ComplexSample)) outputFIFO <- mkSizedBRAMFIFO(1);

  // rule for the first stage
  rule stage1;
    Vector#(TAdd#(1, FFT_LOG_POINTS), Vector#(FFT_POINTS, ComplexSample)) stage_data = newVector();
    stage_data[0] = inputFIFO.first();
    inputFIFO.deq();
    stage_data[1] = stage_f(0, stage_data[0]);
    isb1.enq(stage_data[1]);
  endrule

  rule stage2;
  Vector#(TAdd#(1, FFT_LOG_POINTS), Vector#(FFT_POINTS, ComplexSample)) stage_data = newVector();
  stage_data[1] = isb1.first;
  isb1.deq;
  stage_data[2] = stage_f(1, stage_data[1]);
  isb2.enq(stage_data[2]);
  endrule

  // rule for last stage
  rule stage3;
    Vector#(TAdd#(1, FFT_LOG_POINTS), Vector#(FFT_POINTS, ComplexSample)) stage_data = newVector();
    stage_data[2] = isb2.first;
    isb2.deq;
    stage_data[3] = stage_f(2, stage_data[2]);
    outputFIFO.enq(stage_data[valueof(FFT_LOG_POINTS)]);
  endrule

  interface Put request;
    method Action put(Vector#(FFT_POINTS, ComplexSample) x);
        inputFIFO.enq(bitReverse(x));
    endmethod
  endinterface

  interface Get response = toGet(outputFIFO);

endmodule

module mkAECombinationalFFT (FFT);

  // Statically generate the twiddle factors table.
  TwiddleTable twiddles = genTwiddles();

  // Define the stage_f function which uses the generated twiddles.
  function Vector#(FFT_POINTS, ComplexSample) stage_f(Bit#(TLog#(FFT_LOG_POINTS)) stage, Vector#(FFT_POINTS, ComplexSample) stage_in);
    return ae_stage_ft(twiddles, stage, stage_in);
  endfunction

  FIFO#(Vector#(FFT_POINTS, ComplexSample)) inputFIFO  <- mkSizedBRAMFIFO(1);
  FIFO#(Vector#(FFT_POINTS, ComplexSample)) outputFIFO <- mkSizedBRAMFIFO(1);

  // This rule performs fft using a big mass of combinational logic.
  rule comb_fft;

    Vector#(TAdd#(1, FFT_LOG_POINTS), Vector#(FFT_POINTS, ComplexSample)) stage_data = newVector();
    stage_data[0] = inputFIFO.first();
    inputFIFO.deq();

    // hardcoded for 8-pt fft.
    // for(Integer stage = 0; stage < valueof(FFT_LOG_POINTS); stage=stage+1) begin
    //     stage_data[stage+1] = stage_f(fromInteger(stage), stage_data[stage]);
    // end
    stage_data[1] = stage_f(0, stage_data[0]);
    stage_data[2] = stage_f(1, stage_data[1]);

    outputFIFO.enq(stage_data[valueof(FFT_LOG_POINTS)]);
  endrule

  interface Put request;
    method Action put(Vector#(FFT_POINTS, ComplexSample) x);
        inputFIFO.enq(aebitReverse(x));
    endmethod
  endinterface

  interface Get response = toGet(outputFIFO);

endmodule

// Wrapper around The FFT module we actually want to use
module mkFFT (FFT);
    FFT fft <- mkCombinationalFFT();
    // FFT fft <- mkAECombinationalFFT();
    // FFT fft <- mkPipelinedFFT();

    interface Put request = fft.request;
    interface Get response = fft.response;
endmodule

// Inverse FFT, based on the mkFFT module.
// ifft[k] = fft[N-k]/N
module mkIFFT (FFT);

    FFT fft <- mkFFT();
    FIFO#(Vector#(FFT_POINTS, ComplexSample)) outfifo <- mkSizedBRAMFIFO(1);

    Integer n = valueof(FFT_POINTS);
    Integer lgn = valueof(FFT_LOG_POINTS);

    function ComplexSample scaledown(ComplexSample x);
        return cmplx(x.rel >> lgn, x.img >> lgn);
    endfunction

    rule inversify (True);
        let x <- fft.response.get();
        Vector#(FFT_POINTS, ComplexSample) rx = newVector;

        for (Integer i = 0; i < n; i = i+1) begin
            rx[i] = x[(n - i)%n];
        end
        outfifo.enq(map(scaledown, rx));
    endrule

    interface Put request = fft.request;
    interface Get response = toGet(outfifo);

endmodule

